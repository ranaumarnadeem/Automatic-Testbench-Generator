module priority_encoder_8(
    input [7:0] in,
    input en,
    output reg [2:0] out,
    output reg valid
);
    always @(*) begin
        if (!en) begin
            out = 3'b000;
            valid = 0;
        end else begin
            valid = 1;
            casex (in)
                8'b1xxxxxxx: out = 3'b111;
                8'b01xxxxxx: out = 3'b110;
                8'b001xxxxx: out = 3'b101;
                8'b0001xxxx: out = 3'b100;
                8'b00001xxx: out = 3'b011;
                8'b000001xx: out = 3'b010;
                8'b0000001x: out = 3'b001;
                8'b00000001: out = 3'b000;
                default: begin out = 3'b000; valid = 0; end
            endcase
        end
    end
endmodule



// ---- Auto-generated testbench ----
`timescale 1ns/1ps
module priority_encoder_8_tb;
// Declare inputs and outputs
    reg [7:0] in;
    reg en;
    wire [2:0] out;
    wire valid;

// Instantiate DUT
    priority_encoder_8 uut (
        .in(in),
        .en(en),
        .out(out),
        .valid(valid)
    );

initial begin
        #10 in = 0; en = 0;
        #10 in = 0; en = 1;
        #10 in = 1; en = 0;
        #10 in = 1; en = 1;
        #10 in = 2; en = 0;
        #10 in = 2; en = 1;
        #10 in = 3; en = 0;
        #10 in = 3; en = 1;
        #10 in = 4; en = 0;
        #10 in = 4; en = 1;
        #10 in = 5; en = 0;
        #10 in = 5; en = 1;
        #10 in = 6; en = 0;
        #10 in = 6; en = 1;
        #10 in = 7; en = 0;
        #10 in = 7; en = 1;
        #10 in = 8; en = 0;
        #10 in = 8; en = 1;
        #10 in = 9; en = 0;
        #10 in = 9; en = 1;
        #10 in = 10; en = 0;
        #10 in = 10; en = 1;
        #10 in = 11; en = 0;
        #10 in = 11; en = 1;
        #10 in = 12; en = 0;
        #10 in = 12; en = 1;
        #10 in = 13; en = 0;
        #10 in = 13; en = 1;
        #10 in = 14; en = 0;
        #10 in = 14; en = 1;
        #10 in = 15; en = 0;
        #10 in = 15; en = 1;
        #10 in = 16; en = 0;
        #10 in = 16; en = 1;
        #10 in = 17; en = 0;
        #10 in = 17; en = 1;
        #10 in = 18; en = 0;
        #10 in = 18; en = 1;
        #10 in = 19; en = 0;
        #10 in = 19; en = 1;
        #10 in = 20; en = 0;
        #10 in = 20; en = 1;
        #10 in = 21; en = 0;
        #10 in = 21; en = 1;
        #10 in = 22; en = 0;
        #10 in = 22; en = 1;
        #10 in = 23; en = 0;
        #10 in = 23; en = 1;
        #10 in = 24; en = 0;
        #10 in = 24; en = 1;
        #10 in = 25; en = 0;
        #10 in = 25; en = 1;
        #10 in = 26; en = 0;
        #10 in = 26; en = 1;
        #10 in = 27; en = 0;
        #10 in = 27; en = 1;
        #10 in = 28; en = 0;
        #10 in = 28; en = 1;
        #10 in = 29; en = 0;
        #10 in = 29; en = 1;
        #10 in = 30; en = 0;
        #10 in = 30; en = 1;
        #10 in = 31; en = 0;
        #10 in = 31; en = 1;
        #10 in = 32; en = 0;
        #10 in = 32; en = 1;
        #10 in = 33; en = 0;
        #10 in = 33; en = 1;
        #10 in = 34; en = 0;
        #10 in = 34; en = 1;
        #10 in = 35; en = 0;
        #10 in = 35; en = 1;
        #10 in = 36; en = 0;
        #10 in = 36; en = 1;
        #10 in = 37; en = 0;
        #10 in = 37; en = 1;
        #10 in = 38; en = 0;
        #10 in = 38; en = 1;
        #10 in = 39; en = 0;
        #10 in = 39; en = 1;
        #10 in = 40; en = 0;
        #10 in = 40; en = 1;
        #10 in = 41; en = 0;
        #10 in = 41; en = 1;
        #10 in = 42; en = 0;
        #10 in = 42; en = 1;
        #10 in = 43; en = 0;
        #10 in = 43; en = 1;
        #10 in = 44; en = 0;
        #10 in = 44; en = 1;
        #10 in = 45; en = 0;
        #10 in = 45; en = 1;
        #10 in = 46; en = 0;
        #10 in = 46; en = 1;
        #10 in = 47; en = 0;
        #10 in = 47; en = 1;
        #10 in = 48; en = 0;
        #10 in = 48; en = 1;
        #10 in = 49; en = 0;
        #10 in = 49; en = 1;
        #10 in = 50; en = 0;
        #10 in = 50; en = 1;
        #10 in = 51; en = 0;
        #10 in = 51; en = 1;
        #10 in = 52; en = 0;
        #10 in = 52; en = 1;
        #10 in = 53; en = 0;
        #10 in = 53; en = 1;
        #10 in = 54; en = 0;
        #10 in = 54; en = 1;
        #10 in = 55; en = 0;
        #10 in = 55; en = 1;
        #10 in = 56; en = 0;
        #10 in = 56; en = 1;
        #10 in = 57; en = 0;
        #10 in = 57; en = 1;
        #10 in = 58; en = 0;
        #10 in = 58; en = 1;
        #10 in = 59; en = 0;
        #10 in = 59; en = 1;
        #10 in = 60; en = 0;
        #10 in = 60; en = 1;
        #10 in = 61; en = 0;
        #10 in = 61; en = 1;
        #10 in = 62; en = 0;
        #10 in = 62; en = 1;
        #10 in = 63; en = 0;
        #10 in = 63; en = 1;
        #10 in = 64; en = 0;
        #10 in = 64; en = 1;
        #10 in = 65; en = 0;
        #10 in = 65; en = 1;
        #10 in = 66; en = 0;
        #10 in = 66; en = 1;
        #10 in = 67; en = 0;
        #10 in = 67; en = 1;
        #10 in = 68; en = 0;
        #10 in = 68; en = 1;
        #10 in = 69; en = 0;
        #10 in = 69; en = 1;
        #10 in = 70; en = 0;
        #10 in = 70; en = 1;
        #10 in = 71; en = 0;
        #10 in = 71; en = 1;
        #10 in = 72; en = 0;
        #10 in = 72; en = 1;
        #10 in = 73; en = 0;
        #10 in = 73; en = 1;
        #10 in = 74; en = 0;
        #10 in = 74; en = 1;
        #10 in = 75; en = 0;
        #10 in = 75; en = 1;
        #10 in = 76; en = 0;
        #10 in = 76; en = 1;
        #10 in = 77; en = 0;
        #10 in = 77; en = 1;
        #10 in = 78; en = 0;
        #10 in = 78; en = 1;
        #10 in = 79; en = 0;
        #10 in = 79; en = 1;
        #10 in = 80; en = 0;
        #10 in = 80; en = 1;
        #10 in = 81; en = 0;
        #10 in = 81; en = 1;
        #10 in = 82; en = 0;
        #10 in = 82; en = 1;
        #10 in = 83; en = 0;
        #10 in = 83; en = 1;
        #10 in = 84; en = 0;
        #10 in = 84; en = 1;
        #10 in = 85; en = 0;
        #10 in = 85; en = 1;
        #10 in = 86; en = 0;
        #10 in = 86; en = 1;
        #10 in = 87; en = 0;
        #10 in = 87; en = 1;
        #10 in = 88; en = 0;
        #10 in = 88; en = 1;
        #10 in = 89; en = 0;
        #10 in = 89; en = 1;
        #10 in = 90; en = 0;
        #10 in = 90; en = 1;
        #10 in = 91; en = 0;
        #10 in = 91; en = 1;
        #10 in = 92; en = 0;
        #10 in = 92; en = 1;
        #10 in = 93; en = 0;
        #10 in = 93; en = 1;
        #10 in = 94; en = 0;
        #10 in = 94; en = 1;
        #10 in = 95; en = 0;
        #10 in = 95; en = 1;
        #10 in = 96; en = 0;
        #10 in = 96; en = 1;
        #10 in = 97; en = 0;
        #10 in = 97; en = 1;
        #10 in = 98; en = 0;
        #10 in = 98; en = 1;
        #10 in = 99; en = 0;
        #10 in = 99; en = 1;
        #10 in = 100; en = 0;
        #10 in = 100; en = 1;
        #10 in = 101; en = 0;
        #10 in = 101; en = 1;
        #10 in = 102; en = 0;
        #10 in = 102; en = 1;
        #10 in = 103; en = 0;
        #10 in = 103; en = 1;
        #10 in = 104; en = 0;
        #10 in = 104; en = 1;
        #10 in = 105; en = 0;
        #10 in = 105; en = 1;
        #10 in = 106; en = 0;
        #10 in = 106; en = 1;
        #10 in = 107; en = 0;
        #10 in = 107; en = 1;
        #10 in = 108; en = 0;
        #10 in = 108; en = 1;
        #10 in = 109; en = 0;
        #10 in = 109; en = 1;
        #10 in = 110; en = 0;
        #10 in = 110; en = 1;
        #10 in = 111; en = 0;
        #10 in = 111; en = 1;
        #10 in = 112; en = 0;
        #10 in = 112; en = 1;
        #10 in = 113; en = 0;
        #10 in = 113; en = 1;
        #10 in = 114; en = 0;
        #10 in = 114; en = 1;
        #10 in = 115; en = 0;
        #10 in = 115; en = 1;
        #10 in = 116; en = 0;
        #10 in = 116; en = 1;
        #10 in = 117; en = 0;
        #10 in = 117; en = 1;
        #10 in = 118; en = 0;
        #10 in = 118; en = 1;
        #10 in = 119; en = 0;
        #10 in = 119; en = 1;
        #10 in = 120; en = 0;
        #10 in = 120; en = 1;
        #10 in = 121; en = 0;
        #10 in = 121; en = 1;
        #10 in = 122; en = 0;
        #10 in = 122; en = 1;
        #10 in = 123; en = 0;
        #10 in = 123; en = 1;
        #10 in = 124; en = 0;
        #10 in = 124; en = 1;
        #10 in = 125; en = 0;
        #10 in = 125; en = 1;
        #10 in = 126; en = 0;
        #10 in = 126; en = 1;
        #10 in = 127; en = 0;
        #10 in = 127; en = 1;
        #10 in = 128; en = 0;
        #10 in = 128; en = 1;
        #10 in = 129; en = 0;
        #10 in = 129; en = 1;
        #10 in = 130; en = 0;
        #10 in = 130; en = 1;
        #10 in = 131; en = 0;
        #10 in = 131; en = 1;
        #10 in = 132; en = 0;
        #10 in = 132; en = 1;
        #10 in = 133; en = 0;
        #10 in = 133; en = 1;
        #10 in = 134; en = 0;
        #10 in = 134; en = 1;
        #10 in = 135; en = 0;
        #10 in = 135; en = 1;
        #10 in = 136; en = 0;
        #10 in = 136; en = 1;
        #10 in = 137; en = 0;
        #10 in = 137; en = 1;
        #10 in = 138; en = 0;
        #10 in = 138; en = 1;
        #10 in = 139; en = 0;
        #10 in = 139; en = 1;
        #10 in = 140; en = 0;
        #10 in = 140; en = 1;
        #10 in = 141; en = 0;
        #10 in = 141; en = 1;
        #10 in = 142; en = 0;
        #10 in = 142; en = 1;
        #10 in = 143; en = 0;
        #10 in = 143; en = 1;
        #10 in = 144; en = 0;
        #10 in = 144; en = 1;
        #10 in = 145; en = 0;
        #10 in = 145; en = 1;
        #10 in = 146; en = 0;
        #10 in = 146; en = 1;
        #10 in = 147; en = 0;
        #10 in = 147; en = 1;
        #10 in = 148; en = 0;
        #10 in = 148; en = 1;
        #10 in = 149; en = 0;
        #10 in = 149; en = 1;
        #10 in = 150; en = 0;
        #10 in = 150; en = 1;
        #10 in = 151; en = 0;
        #10 in = 151; en = 1;
        #10 in = 152; en = 0;
        #10 in = 152; en = 1;
        #10 in = 153; en = 0;
        #10 in = 153; en = 1;
        #10 in = 154; en = 0;
        #10 in = 154; en = 1;
        #10 in = 155; en = 0;
        #10 in = 155; en = 1;
        #10 in = 156; en = 0;
        #10 in = 156; en = 1;
        #10 in = 157; en = 0;
        #10 in = 157; en = 1;
        #10 in = 158; en = 0;
        #10 in = 158; en = 1;
        #10 in = 159; en = 0;
        #10 in = 159; en = 1;
        #10 in = 160; en = 0;
        #10 in = 160; en = 1;
        #10 in = 161; en = 0;
        #10 in = 161; en = 1;
        #10 in = 162; en = 0;
        #10 in = 162; en = 1;
        #10 in = 163; en = 0;
        #10 in = 163; en = 1;
        #10 in = 164; en = 0;
        #10 in = 164; en = 1;
        #10 in = 165; en = 0;
        #10 in = 165; en = 1;
        #10 in = 166; en = 0;
        #10 in = 166; en = 1;
        #10 in = 167; en = 0;
        #10 in = 167; en = 1;
        #10 in = 168; en = 0;
        #10 in = 168; en = 1;
        #10 in = 169; en = 0;
        #10 in = 169; en = 1;
        #10 in = 170; en = 0;
        #10 in = 170; en = 1;
        #10 in = 171; en = 0;
        #10 in = 171; en = 1;
        #10 in = 172; en = 0;
        #10 in = 172; en = 1;
        #10 in = 173; en = 0;
        #10 in = 173; en = 1;
        #10 in = 174; en = 0;
        #10 in = 174; en = 1;
        #10 in = 175; en = 0;
        #10 in = 175; en = 1;
        #10 in = 176; en = 0;
        #10 in = 176; en = 1;
        #10 in = 177; en = 0;
        #10 in = 177; en = 1;
        #10 in = 178; en = 0;
        #10 in = 178; en = 1;
        #10 in = 179; en = 0;
        #10 in = 179; en = 1;
        #10 in = 180; en = 0;
        #10 in = 180; en = 1;
        #10 in = 181; en = 0;
        #10 in = 181; en = 1;
        #10 in = 182; en = 0;
        #10 in = 182; en = 1;
        #10 in = 183; en = 0;
        #10 in = 183; en = 1;
        #10 in = 184; en = 0;
        #10 in = 184; en = 1;
        #10 in = 185; en = 0;
        #10 in = 185; en = 1;
        #10 in = 186; en = 0;
        #10 in = 186; en = 1;
        #10 in = 187; en = 0;
        #10 in = 187; en = 1;
        #10 in = 188; en = 0;
        #10 in = 188; en = 1;
        #10 in = 189; en = 0;
        #10 in = 189; en = 1;
        #10 in = 190; en = 0;
        #10 in = 190; en = 1;
        #10 in = 191; en = 0;
        #10 in = 191; en = 1;
        #10 in = 192; en = 0;
        #10 in = 192; en = 1;
        #10 in = 193; en = 0;
        #10 in = 193; en = 1;
        #10 in = 194; en = 0;
        #10 in = 194; en = 1;
        #10 in = 195; en = 0;
        #10 in = 195; en = 1;
        #10 in = 196; en = 0;
        #10 in = 196; en = 1;
        #10 in = 197; en = 0;
        #10 in = 197; en = 1;
        #10 in = 198; en = 0;
        #10 in = 198; en = 1;
        #10 in = 199; en = 0;
        #10 in = 199; en = 1;
        #10 in = 200; en = 0;
        #10 in = 200; en = 1;
        #10 in = 201; en = 0;
        #10 in = 201; en = 1;
        #10 in = 202; en = 0;
        #10 in = 202; en = 1;
        #10 in = 203; en = 0;
        #10 in = 203; en = 1;
        #10 in = 204; en = 0;
        #10 in = 204; en = 1;
        #10 in = 205; en = 0;
        #10 in = 205; en = 1;
        #10 in = 206; en = 0;
        #10 in = 206; en = 1;
        #10 in = 207; en = 0;
        #10 in = 207; en = 1;
        #10 in = 208; en = 0;
        #10 in = 208; en = 1;
        #10 in = 209; en = 0;
        #10 in = 209; en = 1;
        #10 in = 210; en = 0;
        #10 in = 210; en = 1;
        #10 in = 211; en = 0;
        #10 in = 211; en = 1;
        #10 in = 212; en = 0;
        #10 in = 212; en = 1;
        #10 in = 213; en = 0;
        #10 in = 213; en = 1;
        #10 in = 214; en = 0;
        #10 in = 214; en = 1;
        #10 in = 215; en = 0;
        #10 in = 215; en = 1;
        #10 in = 216; en = 0;
        #10 in = 216; en = 1;
        #10 in = 217; en = 0;
        #10 in = 217; en = 1;
        #10 in = 218; en = 0;
        #10 in = 218; en = 1;
        #10 in = 219; en = 0;
        #10 in = 219; en = 1;
        #10 in = 220; en = 0;
        #10 in = 220; en = 1;
        #10 in = 221; en = 0;
        #10 in = 221; en = 1;
        #10 in = 222; en = 0;
        #10 in = 222; en = 1;
        #10 in = 223; en = 0;
        #10 in = 223; en = 1;
        #10 in = 224; en = 0;
        #10 in = 224; en = 1;
        #10 in = 225; en = 0;
        #10 in = 225; en = 1;
        #10 in = 226; en = 0;
        #10 in = 226; en = 1;
        #10 in = 227; en = 0;
        #10 in = 227; en = 1;
        #10 in = 228; en = 0;
        #10 in = 228; en = 1;
        #10 in = 229; en = 0;
        #10 in = 229; en = 1;
        #10 in = 230; en = 0;
        #10 in = 230; en = 1;
        #10 in = 231; en = 0;
        #10 in = 231; en = 1;
        #10 in = 232; en = 0;
        #10 in = 232; en = 1;
        #10 in = 233; en = 0;
        #10 in = 233; en = 1;
        #10 in = 234; en = 0;
        #10 in = 234; en = 1;
        #10 in = 235; en = 0;
        #10 in = 235; en = 1;
        #10 in = 236; en = 0;
        #10 in = 236; en = 1;
        #10 in = 237; en = 0;
        #10 in = 237; en = 1;
        #10 in = 238; en = 0;
        #10 in = 238; en = 1;
        #10 in = 239; en = 0;
        #10 in = 239; en = 1;
        #10 in = 240; en = 0;
        #10 in = 240; en = 1;
        #10 in = 241; en = 0;
        #10 in = 241; en = 1;
        #10 in = 242; en = 0;
        #10 in = 242; en = 1;
        #10 in = 243; en = 0;
        #10 in = 243; en = 1;
        #10 in = 244; en = 0;
        #10 in = 244; en = 1;
        #10 in = 245; en = 0;
        #10 in = 245; en = 1;
        #10 in = 246; en = 0;
        #10 in = 246; en = 1;
        #10 in = 247; en = 0;
        #10 in = 247; en = 1;
        #10 in = 248; en = 0;
        #10 in = 248; en = 1;
        #10 in = 249; en = 0;
        #10 in = 249; en = 1;
        #10 in = 250; en = 0;
        #10 in = 250; en = 1;
        #10 in = 251; en = 0;
        #10 in = 251; en = 1;
        #10 in = 252; en = 0;
        #10 in = 252; en = 1;
        #10 in = 253; en = 0;
        #10 in = 253; en = 1;
        #10 in = 254; en = 0;
        #10 in = 254; en = 1;
        #10 in = 255; en = 0;
        #10 in = 255; en = 1;
        $finish;
end
endmodule